LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY LAST_XOR IS PORT
(
V0_IN :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
V1_IN :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
V2_IN :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
V3_IN :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
HASH :OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
);
END LAST_XOR;
ARCHITECTURE ARCH_LAST_XOR OF LAST_XOR IS
BEGIN
HASH <= V0_IN XOR V1_IN XOR V2_IN XOR V3_IN;
END ARCHITECTURE;