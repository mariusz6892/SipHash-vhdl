LIBRARY IEEE  ; 
LIBRARY STD   ; 
LIBRARY WORK  ; 
USE IEEE.NUMERIC_STD.ALL  ; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_TEXTIO.ALL  ; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL  ; 
USE STD.TEXTIO.ALL  ; 
USE WORK.ALL  ; 
ENTITY SIPROUND_TB  IS 
END ; 
 
ARCHITECTURE SIPROUND_TB_ARCH OF SIPROUND_TB IS
	SIGNAL V0_IN : STD_LOGIC_VECTOR(63 DOWNTO 0); 
	SIGNAL V1_IN :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL V2_IN :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL V3_IN :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL V0_OUT :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL V1_OUT  :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL V2_OUT  :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL V3_OUT  :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL CLKp :time := 40 ns;
	SIGNAL clk :STD_LOGIC;
	
	COMPONENT SIPROUND IS PORT
(	
	V0_IN :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
	V1_IN :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
	V2_IN :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
	V3_IN :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
	V0_OUT :OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
	V1_OUT :OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
	V2_OUT :OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
	V3_OUT :OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	DUT : SIPROUND  
	PORT MAP 
	( 
		V0_IN   => V0_IN,		
		V1_IN => V1_IN,
		V2_IN => V2_IN,
		V3_IN => V3_IN,
		V0_OUT => V0_OUT,
		V1_OUT => V1_OUT,
		V2_OUT => V2_OUT,
		V3_OUT => V3_OUT
	); 
	
	Process
	Begin
		clk  <= '0'  ; wait for CLKp/2;
		clk  <= '1'  ; wait for CLKp/2;
	End Process;
	
	PROCESS
	BEGIN
	V0_IN <= X"FFFFFFFFFFFFFFFF"; V1_IN <= X"1111111111111111"; V2_IN <= X"FFFFFFFFFFFFFFFF"; V3_IN <= X"1111111111111111"; wait for CLKp;
	V0_IN <= X"FFFFA02301010230"; V1_IN <= X"12341AD4123456AD"; V2_IN <= X"BCD232543141123A"; V3_IN <= X"FEAD234131231ADE"; wait for CLKp;
	END PROCESS;
	

END;
