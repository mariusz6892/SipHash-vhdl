LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY SIPHASH IS PORT
(
MESSAGE_0 :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
MESSAGE_1 :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
KEY_0 :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
KEY_1 :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
HASH :OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
);
END SIPHASH;
ARCHITECTURE ARCH_SIPHASH OF SIPHASH IS
SIGNAL V_0 :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_1 :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_2 :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_3 :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_0_AFTER1SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_1_AFTER1SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_2_AFTER1SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_3_AFTER1SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_0_AFTER2SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_1_AFTER2SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_2_AFTER2SR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_3_AFTER2SR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_0_AFTERMXOR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_3_AFTERMXOR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_0_AFTER3SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_1_AFTER3SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_2_AFTER3SR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_3_AFTER3SR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_0_AFTER4SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_1_AFTER4SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_2_AFTER4SR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_3_AFTER4SR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_0_AFTERLMXOR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_2_AFTERLMXOR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_0_AFTER5SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_1_AFTER5SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_2_AFTER5SR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_3_AFTER5SR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_0_AFTER6SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_1_AFTER6SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_2_AFTER6SR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_3_AFTER6SR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_0_AFTER7SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_1_AFTER7SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_2_AFTER7SR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_3_AFTER7SR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_0_AFTER8SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_1_AFTER8SR :STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_2_AFTER8SR:STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL V_3_AFTER8SR:STD_LOGIC_VECTOR(63 DOWNTO 0);

BEGIN
INITIAL_XOR			: ENTITY WORK.INITIAL_XOR 			PORT MAP(KEY_0,KEY_1,MESSAGE_0,V_0,V_1,V_2,V_3);
SIPROUND_1 			: ENTITY WORK.SIPROUND    			PORT MAP(V_0,V_1,V_2,V_3,V_0_AFTER1SR,V_1_AFTER1SR,V_2_AFTER1SR,V_3_AFTER1SR);
SIPROUND_2			: ENTITY WORK.SIPROUND	 			PORT MAP(V_0_AFTER1SR,V_1_AFTER1SR,V_2_AFTER1SR,V_3_AFTER1SR,V_0_AFTER2SR,V_1_AFTER2SR,V_2_AFTER2SR,V_3_AFTER2SR);
MIDDLE_XOR 			: ENTITY WORK.MIDDLE_XOR 			PORT MAP(V_0_AFTER2SR,V_3_AFTER2SR,MESSAGE_0,MESSAGE_1,V_0_AFTERMXOR,V_3_AFTERMXOR);
SIPROUND_3 			: ENTITY WORK.SIPROUND   			PORT MAP(V_0_AFTERMXOR,V_1_AFTER2SR,V_2_AFTER2SR,V_3_AFTERMXOR,V_0_AFTER3SR,V_1_AFTER3SR,V_2_AFTER3SR,V_3_AFTER3SR);
SIPROUND_4 			: ENTITY WORK.SIPROUND    			PORT MAP(V_0_AFTER3SR,V_1_AFTER3SR,V_2_AFTER3SR,V_3_AFTER3SR,V_0_AFTER4SR,V_1_AFTER4SR,V_2_AFTER4SR,V_3_AFTER4SR);
LASTMESSAGE_XOR   : ENTITY WORK.LASTMESSAGE_XOR  	PORT MAP(V_0_AFTER4SR,V_2_AFTER4SR,MESSAGE_1,V_0_AFTERLMXOR,V_2_AFTERLMXOR);
SIPROUND_5 			: ENTITY WORK.SIPROUND   			PORT MAP(V_0_AFTERLMXOR,V_1_AFTER4SR,V_2_AFTERLMXOR,V_3_AFTER4SR,V_0_AFTER5SR,V_1_AFTER5SR,V_2_AFTER5SR,V_3_AFTER5SR);
SIPROUND_6 			: ENTITY WORK.SIPROUND   			PORT MAP(V_0_AFTER5SR,V_1_AFTER5SR,V_2_AFTER5SR,V_3_AFTER5SR,V_0_AFTER6SR,V_1_AFTER6SR,V_2_AFTER6SR,V_3_AFTER6SR);
SIPROUND_7 			: ENTITY WORK.SIPROUND   			PORT MAP(V_0_AFTER6SR,V_1_AFTER6SR,V_2_AFTER6SR,V_3_AFTER6SR,V_0_AFTER7SR,V_1_AFTER7SR,V_2_AFTER7SR,V_3_AFTER7SR);
SIPROUND_8 			: ENTITY WORK.SIPROUND   			PORT MAP(V_0_AFTER7SR,V_1_AFTER7SR,V_2_AFTER7SR,V_3_AFTER7SR,V_0_AFTER8SR,V_1_AFTER8SR,V_2_AFTER8SR,V_3_AFTER8SR);
LAST_XOR				: ENTITY WORK.LAST_XOR				PORT MAP(V_0_AFTER8SR,V_1_AFTER8SR,V_2_AFTER8SR,V_3_AFTER8SR,HASH);
END ARCHITECTURE;