----------------------------------
-- Łukasz DZIEŁ (883533374)     --
-- FPGACOMMEXAMPLE-v2           --
-- 01.2016                      --
-- 1.0                          --
----------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY WORK;
USE WORK.ALL;

ENTITY FPGAX IS PORT
(	
	CLK				:IN STD_LOGIC;
	RS232_TX			:OUT STD_LOGIC;
	RS232_RX			:IN STD_LOGIC); END ENTITY;


ARCHITECTURE FPGAX_ARCH OF FPGAX IS	
	
	SIGNAL ZERO :STD_LOGIC; 
	
	SIGNAL TEMP1 :STD_LOGIC;
	SIGNAL TEMP2 :STD_LOGIC;
	
	SIGNAL TEMP3 :STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL TEMP4 :STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL TEMP5 :STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	SIGNAL NRBYTES 	:STD_LOGIC_VECTOR(3  DOWNTO 0);
	SIGNAL MESSAGE 	:STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL KEY_0		:STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL KEY_1		:STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL HASH			:STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL HASH_READY	:STD_LOGIC;
	
BEGIN
	ZERO <= '0';
	
	unit00: ENTITY WORK.RS232_STANDARD_INTERFACE PORT MAP (
			CLK		=> CLK,
			INIT		=> ZERO,
			TX			=> RS232_TX,
			RX			=> RS232_RX,
			INT_WR	=> TEMP1,
			INT_RD	=> TEMP2,
			INT_ADDR	=> TEMP3,
			INT_DIN	=> TEMP4,
			INT_DOUT	=> TEMP5);
	
	example01: ENTITY WORK.EXAMPLEX PORT MAP (
			CLK	=> CLK,
			INIT	=> ZERO,
			RD		=> TEMP2,
			WR		=> TEMP1,
			ADDR	=> TEMP3,
			DIN	=> TEMP5,
			DOUT	=> TEMP4,
			NRBYTES 		=> NRBYTES,
			MESSAGE 		=> MESSAGE,
			KEY_0	  		=> KEY_0,
			KEY_1   		=> KEY_1,
			HASH   		=> HASH,
			HASH_READY  => HASH_READY);
			
	siphashstates02: ENTITY WORK.SIPHASHSTATES PORT MAP (
			CLK 			=> CLK,
			MESSAGE 		=> MESSAGE,
			KEY_0	  		=> KEY_0,
			KEY_1   		=> KEY_1,
			NRBYTES 		=> NRBYTES,
			HASH   		=> HASH,
			HASH_READY  => HASH_READY);
	
END ARCHITECTURE;