LIBRARY IEEE  ; 
LIBRARY STD   ; 
LIBRARY WORK  ; 
USE IEEE.NUMERIC_STD.ALL  ; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_TEXTIO.ALL  ; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL  ; 
USE STD.TEXTIO.ALL  ; 
USE WORK.ALL  ; 
ENTITY EXAMPLE2_TB  IS 
END ; 
 
ARCHITECTURE EXAMPLE2_TB_ATCH OF EXAMPLE2_TB IS
	SIGNAL WR : STD_LOGIC; 
	SIGNAL INIT: STD_LOGIC;
	SIGNAL CLK : STD_LOGIC; 
	SIGNAL RD : STD_LOGIC; 
	SIGNAL ADDR : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL DIN : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL DOUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL NRBYTES :STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL MESSAGE :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL KEY_0 :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL KEY_1 :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL HASH  :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL HASH_READY :STD_LOGIC;
	
	SIGNAL CLKp : time:=40ns;
	
	COMPONENT EXAMPLEX IS PORT
(	
	CLK	:IN STD_LOGIC;
	INIT	:IN STD_LOGIC;
	RD   	:IN STD_LOGIC;
	WR		:IN STD_LOGIC;
	ADDR	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DIN	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DOUT	:OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	NRBYTES 		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	MESSAGE 		: OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
	KEY_0	  		: OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
	KEY_1   		: OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
	
	HASH   		: IN STD_LOGIC_VECTOR(63 DOWNTO 0);
	HASH_READY  : IN STD_LOGIC
	);
	END COMPONENT;

BEGIN
	DUT : EXAMPLEX  
	PORT MAP 
	( 
		CLK   => CLK,
		INIT  => INIT,
		WR => WR,
		RD => RD,
		ADDR => ADDR,
		DIN => DIN,
		DOUT => DOUT,
		
		NRBYTES => NRBYTES,
		MESSAGE => MESSAGE,
		KEY_0 => KEY_0,
		KEY_1 => KEY_1,
		HASH => HASH,
		HASH_READY => HASH_READY
	); 

	Process
	Begin
		clk  <= '0'  ; wait for CLKp/2;
		clk  <= '1'  ; wait for CLKp/2;
	End Process;
	
	PROCESS
	BEGIN
	WR <= '1'; ADDR <= X"00000000"; DIN <= X"00000008"; wait for CLKp;
	WR <= '1'; ADDR <= X"00000001"; DIN <= X"6b6f6c61"; wait for CLKp;
	WR <= '1'; ADDR <= X"00000002"; DIN <= X"626f7261"; wait for CLKp;
	WR <= '1'; ADDR <= X"00000003"; DIN <= X"636a616d"; wait for CLKp;
	WR <= '1'; ADDR <= X"00000004"; DIN <= X"616d6178"; wait for CLKp;
	WR <= '1'; ADDR <= X"00000005"; DIN <= X"68656c6c"; wait for CLKp;
	WR <= '1'; ADDR <= X"00000006"; DIN <= X"6f6d616d"; wait for CLKp;
	WR <= '0'; wait for CLKp;
	
	HASH_READY <='1'; HASH <= X"0123456789ABCDEF"; wait for CLKp;
	
	RD <= '1'; ADDR <= X"00000007";wait for CLKp;
	RD <= '0'; wait for CLKp;
	RD <= '1'; ADDR <= X"00000008";wait for CLKp;
	RD <= '0'; wait for CLKp;
	
	WAIT;
	END PROCESS;
	

END;
