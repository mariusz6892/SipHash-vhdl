----------------------------------
-- Łukasz DZIEŁ (883533374)     --
-- FPGACOMMEXAMPLE-v2           --
-- 01.2016                      --
-- 1.0                          --
----------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY EXAMPLE IS PORT
(	
	CLK	:IN STD_LOGIC;
	INIT	:IN STD_LOGIC;
	RD   	:IN STD_LOGIC;
	WR		:IN STD_LOGIC;
	ADDR	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DIN	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DOUT	:OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	
);
END ENTITY;

ARCHITECTURE EXAMPLE_ARCH OF EXAMPLE IS
	
	TYPE MEMORY_BLOCK IS ARRAY (0 TO 15) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MEM : MEMORY_BLOCK;
	
	SIGNAL MESSAGE_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
	SIGNAL MESSAGE_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
	SIGNAL KEY_0	  : STD_LOGIC_VECTOR (63 DOWNTO 0);
	SIGNAL KEY_1     : STD_LOGIC_VECTOR (63 DOWNTO 0);
	SIGNAL HASH      : STD_LOGIC_VECTOR (63 DOWNTO 0);
	
BEGIN
	
	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF (WR = '1') THEN
				MEM(conv_integer(ADDR)) <= DIN;
			ELSE
				MESSAGE_0 <=MEM(conv_integer(X"00000000")) & MEM(conv_integer(X"00000001"));
				MESSAGE_1 <=MEM(conv_integer(X"00000002")) & MEM(conv_integer(X"00000003"));
				KEY_0 <=MEM(conv_integer(X"00000004")) & MEM(conv_integer(X"00000005"));
				KEY_1 <=MEM(conv_integer(X"00000006")) & MEM(conv_integer(X"00000007"));
				MEM(conv_integer(X"00000008")) <= HASH(63 DOWNTO 32);
				MEM(conv_integer(X"00000009")) <= HASH(31 DOWNTO 0);
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF(RD = '1') THEN
				DOUT <= MEM(conv_integer(ADDR));
			ELSE
				DOUT <= (others => 'Z');
			END IF;
		END IF;
	END PROCESS;
	
	SIPHASH: ENTITY WORK.SIPHASH PORT MAP(MESSAGE_0, MESSAGE_1, KEY_0, KEY_1, HASH);
	
	
END ARCHITECTURE;