LIBRARY IEEE  ; 
LIBRARY STD   ; 
LIBRARY WORK  ; 
USE IEEE.NUMERIC_STD.ALL  ; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_TEXTIO.ALL  ; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL  ; 
USE STD.TEXTIO.ALL  ; 
USE WORK.ALL  ; 
ENTITY SIPHASHSTATES_TB  IS 
END ; 
 
ARCHITECTURE SIPHASHSTATES_TB_ATCH OF SIPHASHSTATES_TB IS
	SIGNAL CLK : STD_LOGIC; 
	SIGNAL NRBYTES :STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL MESSAGE :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL KEY_0 :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL KEY_1 :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL HASH  :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL HASH_READY :STD_LOGIC;
	
	SIGNAL CLKp : time:=40ns;
	
	COMPONENT SIPHASHSTATES IS PORT
(	
	CLK     :  IN  STD_LOGIC;
	MESSAGE :  IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
	KEY_0   :  IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
	KEY_1   :  IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
	NRBYTES :  IN  STD_LOGIC_VECTOR(3  DOWNTO 0);
				
		
	HASH    		:  OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
	HASH_READY  :  OUT STD_LOGIC
	);
	END COMPONENT;

BEGIN
	DUT : SIPHASHSTATES  
	PORT MAP 
	( 
		CLK   => CLK,		
		NRBYTES => NRBYTES,
		MESSAGE => MESSAGE,
		KEY_0 => KEY_0,
		KEY_1 => KEY_1,
		HASH => HASH,
		HASH_READY => HASH_READY
	); 

	Process
	Begin
		clk  <= '0'  ; wait for CLKp/2;
		clk  <= '1'  ; wait for CLKp/2;
	End Process;
	
	PROCESS
	BEGIN
	MESSAGE <= X"68656c6c6f6d616d"; NRBYTES <= X"8"; KEY_0 <= X"6b6f6c61626f7261"; KEY_1 <= X"636a616d616d6178"; wait for CLKp;
	MESSAGE <= X"00656c6c6f6d616d"; NRBYTES <= X"7"; KEY_0 <= X"6b6f6c61626f7261"; KEY_1 <= X"636a616d616d6178"; wait for CLKp;
	WAIT;
	END PROCESS;
	

END;
