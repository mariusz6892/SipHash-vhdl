----------------------------------
-- Łukasz DZIEŁ (883533374)     --
-- FPGACOMMEXAMPLE-v2           --
-- 01.2016                      --
-- 1.0                          --
----------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY EXAMPLEX IS PORT
(	
	CLK	:IN STD_LOGIC;
	INIT	:IN STD_LOGIC;
	RD   	:IN STD_LOGIC;
	WR		:IN STD_LOGIC;
	ADDR	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DIN	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DOUT	:OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	NRBYTES 		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	MESSAGE 		: OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
	KEY_0	  		: OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
	KEY_1   		: OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
	
	HASH   		: IN STD_LOGIC_VECTOR(63 DOWNTO 0);
	HASH_READY  : IN STD_LOGIC
	
);
END ENTITY;

ARCHITECTURE EXAMPLEX_ARCH OF EXAMPLEX IS
	
	TYPE MEMORY_BLOCK IS ARRAY (0 TO 15) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MEM : MEMORY_BLOCK;
	SIGNAL NRBYT : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL HASHJAZDA : STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL HASHJAZDA2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
	

	
BEGIN	

	HASHJAZDA <= HASH(63 DOWNTO 32);
	HASHJAZDA2 <= HASH(31 DOWNTO 0);
	
	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF (WR = '1') THEN
				MEM(conv_integer(ADDR)) <= DIN;
			--ELSIF (HASH_READY = '1') THEN
			--	MEM(conv_integer(X"00000007")) <= HASH(63 DOWNTO 32);
			--	MEM(conv_integer(X"00000008")) <= HASH(31 DOWNTO 0);
			ELSE
				NRBYT <= MEM(conv_integer(X"00000000"));
				NRBYTES <= NRBYT(3 DOWNTO 0);
				KEY_0   <= MEM(conv_integer(X"00000001")) & MEM(conv_integer(X"00000002"));
				KEY_1   <= MEM(conv_integer(X"00000003")) & MEM(conv_integer(X"00000004"));
				MESSAGE <= MEM(conv_integer(X"00000005")) & MEM(conv_integer(X"00000006"));
				MEM(conv_integer(X"00000007")) <= HASHJAZDA;
				MEM(conv_integer(X"00000008")) <= HASHJAZDA2;
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF(RD = '1') THEN
				DOUT <= MEM(conv_integer(ADDR));
			ELSE
				DOUT <= (others => 'Z');
			END IF;
		END IF;
	END PROCESS;
	
	--SIPHASH: ENTITY WORK.SIPHASH PORT MAP(MESSAGE_0, MESSAGE_1, KEY_0, KEY_1, HASH);
	
	
END ARCHITECTURE;