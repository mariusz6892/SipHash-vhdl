LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY SIPROUND IS PORT
(
V0_IN :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
V1_IN :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
V2_IN :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
V3_IN :IN STD_LOGIC_VECTOR (63 DOWNTO 0);
V0_OUT :OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
V1_OUT :OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
V2_OUT :OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
V3_OUT :OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
);
END SIPROUND;
ARCHITECTURE ARCH_SIPROUND OF SIPROUND IS
BEGIN
  PROCESS(V0_IN, V1_IN, V2_IN, V3_IN)
     VARIABLE V0, V1, V2, V3 : UNSIGNED(63 downto 0);
  begin
    V0 := UNSIGNED(V0_IN);
    V1 := UNSIGNED(V1_IN);
    V2 := UNSIGNED(V2_IN);
    V3 := UNSIGNED(V3_IN);

    V0 := V0 + V1;
    V2 := V2 + V3;
    V1 := ROTATE_LEFT(V1, 13);
    V3 := ROTATE_LEFT(V3, 16);

    V1 := V1 XOR V0;
    V3 := V3 XOR V2;
    V0 := ROTATE_LEFT(V0, 32);

    V0 := V0 + V3;
    V2 := V2 + V1;
    V1 := ROTATE_LEFT(V1, 17);
    V3 := ROTATE_LEFT(V3, 21);

    V1 := V1 XOR V2;
    V3 := V3 XOR V0;
    V2 := ROTATE_LEFT(V2, 32);

    V0_OUT <= STD_LOGIC_VECTOR(V0);
    V1_OUT <= STD_LOGIC_VECTOR(V1);
    V2_OUT <= STD_LOGIC_VECTOR(V2);
    V3_OUT <= STD_LOGIC_VECTOR(V3);
  end process;
END ARCHITECTURE;